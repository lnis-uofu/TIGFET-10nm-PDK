
***************************************
.SUBCKT TIGFET_PCELL_SP15CP15_N1 d pgs g pgd s
.ENDS
