* SPICE NETLIST
***************************************

.SUBCKT tigfet1 d pgs g pgd s
.ENDS
***************************************
.SUBCKT test_cell
** N=1 EP=0 IP=0 FDC=0
** WARNING: BAD DEVICE on layer tgate at location (-2.168,-5.082) in cell test_cell (see extraction report).
*.CALIBRE WARNING BADDEV BAD DEVICE(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
