* SPICE NETLIST
***************************************

.SUBCKT tigfet1 d pgd cg pgs s
.ENDS
***************************************
.SUBCKT TIGFET_PCELL_SP15CP15_N2 D S PGD CG PGS
** N=5 EP=5 IP=0 FDC=1
X0 D PGD CG PGS S tigfet1 $X=42 $Y=13 $D=0
.ENDS
***************************************
.SUBCKT G5_XNOR3_N2 Vdd C Vss A B Z
** N=9 EP=6 IP=50 FDC=10
X0 4 Vdd Vss C Vss TIGFET_PCELL_SP15CP15_N2 $T=180 61 1 180 $X=0 $Y=64
X1 4 Vss Vdd C Vdd TIGFET_PCELL_SP15CP15_N2 $T=124 61 0 0 $X=138 $Y=64
X2 6 Vss Vdd B Vdd TIGFET_PCELL_SP15CP15_N2 $T=456 61 1 180 $X=276 $Y=64
X3 7 Vdd Vss A Vss TIGFET_PCELL_SP15CP15_N2 $T=456 325 1 180 $X=276 $Y=328
X4 6 Vdd Vss B Vss TIGFET_PCELL_SP15CP15_N2 $T=400 61 0 0 $X=414 $Y=64
X5 7 Vss Vdd A Vdd TIGFET_PCELL_SP15CP15_N2 $T=400 325 0 0 $X=414 $Y=328
X6 Z C 7 B 7 TIGFET_PCELL_SP15CP15_N2 $T=870 61 1 180 $X=690 $Y=64
X7 Z 4 7 6 7 TIGFET_PCELL_SP15CP15_N2 $T=870 325 1 180 $X=690 $Y=328
X8 Z C A 6 A TIGFET_PCELL_SP15CP15_N2 $T=814 61 0 0 $X=828 $Y=64
X9 Z 4 A B A TIGFET_PCELL_SP15CP15_N2 $T=814 325 0 0 $X=828 $Y=328
.ENDS
***************************************
