* SPICE NETLIST
***************************************

.SUBCKT tigfet1 d pgd cg pgs s
.ENDS
***************************************
.SUBCKT TIGFET_PCELL_SP15CP15_N3 D S PGD CG PGS
** N=5 EP=5 IP=0 FDC=1
X0 D PGD CG PGS S tigfet1 $X=29 $Y=11 $D=0
.ENDS
***************************************
.SUBCKT G4_MAJ3_N3 Vdd Vss A B C Z
** N=8 EP=6 IP=40 FDC=8
X0 4 Vdd Vss B Vss TIGFET_PCELL_SP15CP15_N3 $T=167 63 1 180 $X=0 $Y=64
X1 5 Vdd Vss A Vss TIGFET_PCELL_SP15CP15_N3 $T=167 371 1 180 $X=0 $Y=372
X2 4 Vss Vdd B Vdd TIGFET_PCELL_SP15CP15_N3 $T=137 63 0 0 $X=138 $Y=64
X3 5 Vss Vdd A Vdd TIGFET_PCELL_SP15CP15_N3 $T=137 371 0 0 $X=138 $Y=372
X4 Z A 5 4 5 TIGFET_PCELL_SP15CP15_N3 $T=581 63 1 180 $X=414 $Y=64
X5 Z C 5 B 5 TIGFET_PCELL_SP15CP15_N3 $T=581 371 1 180 $X=414 $Y=372
X6 Z A A B A TIGFET_PCELL_SP15CP15_N3 $T=551 63 0 0 $X=552 $Y=64
X7 Z C A 4 A TIGFET_PCELL_SP15CP15_N3 $T=551 371 0 0 $X=552 $Y=372
.ENDS
***************************************
