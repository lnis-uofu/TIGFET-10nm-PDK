.SUBCKT TIGFET_PCELL_SP15CP15_N1 d pgd cg pgs s
.ENDS