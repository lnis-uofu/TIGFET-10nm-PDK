* SPICE NETLIST
***************************************

.SUBCKT tigfet1 d pgd cg pgs s
.ENDS
***************************************
.SUBCKT TIGFET_PCELL_SP15CP15_N2 D S PGD CG PGS
** N=5 EP=5 IP=0 FDC=1
X0 D PGD CG PGS S tigfet1 $X=42 $Y=13 $D=0
.ENDS
***************************************
.SUBCKT G4_MAJ3_N2 Vdd Vss A B C Z
** N=8 EP=6 IP=40 FDC=8
X0 4 Vdd Vss B Vss TIGFET_PCELL_SP15CP15_N2 $T=180 61 1 180 $X=0 $Y=64
X1 5 Vdd Vss A Vss TIGFET_PCELL_SP15CP15_N2 $T=180 325 1 180 $X=0 $Y=328
X2 4 Vss Vdd B Vdd TIGFET_PCELL_SP15CP15_N2 $T=124 61 0 0 $X=138 $Y=64
X3 5 Vss Vdd A Vdd TIGFET_PCELL_SP15CP15_N2 $T=124 325 0 0 $X=138 $Y=328
X4 Z A 5 4 5 TIGFET_PCELL_SP15CP15_N2 $T=594 61 1 180 $X=414 $Y=64
X5 Z C 5 B 5 TIGFET_PCELL_SP15CP15_N2 $T=594 325 1 180 $X=414 $Y=328
X6 Z A A B A TIGFET_PCELL_SP15CP15_N2 $T=538 61 0 0 $X=552 $Y=64
X7 Z C A 4 A TIGFET_PCELL_SP15CP15_N2 $T=538 325 0 0 $X=552 $Y=328
.ENDS
***************************************
