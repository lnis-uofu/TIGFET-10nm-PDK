* SPICE NETLIST
***************************************

.SUBCKT tigfet1 d pgd cg pgs s
.ENDS
***************************************
.SUBCKT TIGFET_PCELL_SP15CP15_N1 D S PGD CG PGS
** N=5 EP=5 IP=0 FDC=1
X0 D PGD CG PGS S tigfet1 $X=142 $Y=62 $D=0
.ENDS
***************************************
.SUBCKT G4_XOR2_N1 Vss Vdd A B Z
** N=7 EP=5 IP=40 FDC=8
X0 4 Vss Vdd B Vdd TIGFET_PCELL_SP15CP15_N1 $T=280 172 0 180 $X=0 $Y=64
X1 5 Vdd Vss A Vss TIGFET_PCELL_SP15CP15_N1 $T=280 223 1 180 $X=0 $Y=263
X2 4 Vdd Vss B Vss TIGFET_PCELL_SP15CP15_N1 $T=24 172 1 0 $X=138 $Y=64
X3 5 Vss Vdd A Vdd TIGFET_PCELL_SP15CP15_N1 $T=24 223 0 0 $X=138 $Y=263
X4 Z Vdd B 5 B TIGFET_PCELL_SP15CP15_N1 $T=556 24 1 180 $X=276 $Y=64
X5 Z Vss A B A TIGFET_PCELL_SP15CP15_N1 $T=556 371 0 180 $X=276 $Y=263
X6 Z Vdd 4 A 4 TIGFET_PCELL_SP15CP15_N1 $T=300 24 0 0 $X=414 $Y=64
X7 Z Vss 5 4 5 TIGFET_PCELL_SP15CP15_N1 $T=300 371 1 0 $X=414 $Y=263
.ENDS
***************************************
