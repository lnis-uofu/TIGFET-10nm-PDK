.SUBCKT tigfet1 d pgs g pgd s
.ENDS
***************************************
.SUBCKT TIGFET_PCELL_SP15CP15_N1 1 2 3 4 5 
X0 1 3 4 5 2 tigfet1 
.ENDS
