* SPICE NETLIST
***************************************

.SUBCKT tigfet1 d pgs g pgd s
.ENDS
***************************************
.SUBCKT TEST
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
